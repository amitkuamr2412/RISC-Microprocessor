# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:35 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 03:18:35 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:36 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 03:18:36 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:36 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 03:18:36 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:36 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 03:18:36 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:36 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 03:18:36 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 03:18:36 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 03:18:36 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:01
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:11 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 01:33:11 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:11 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 01:33:11 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
vsim work.toplevel
# vsim work.toplevel 
# Start time: 03:18:50 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# vsim work.toplevel 
# Start time: 02:21:38 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# vsim work.toplevel 
# Start time: 01:33:56 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# vsim work.toplevel 
# Start time: 01:18:02 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
add wave -position insertpoint  \
sim:/toplevel/FSM_control/ir_data \
sim:/toplevel/FSM_control/next_state \
sim:/toplevel/FSM_control/state
add wave -position insertpoint  \
sim:/toplevel/Datapat/memory_block/memory_block
add wave -position insertpoint  \
sim:/toplevel/Datapat/reg_file_block/registers
add wave -position insertpoint  \
sim:/toplevel/clock \
sim:/toplevel/reset
force -freeze sim:/toplevel/clock 1 0, 0 {50 ps} -r 100
force -freeze sim:/toplevel/reset 1 0
run
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
force -freeze sim:/toplevel/reset 0 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(0) 0110000010000001 0
force -freeze sim:/toplevel/Datapat/reg_file_block/registers(0) 0000000000000100 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(4) 0000000000000001 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(5) 0000000000000111 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(0) 0110000001000001 0
add wave -position insertpoint  \
sim:/toplevel/Datapat/t4_block/din \
sim:/toplevel/Datapat/t4_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/t2_block/din \
sim:/toplevel/Datapat/t2_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/t5_block/din \
sim:/toplevel/Datapat/t5_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/xorblock/dout \
sim:/toplevel/Datapat/xorblock/xor_a \
sim:/toplevel/Datapat/xorblock/xor_b
add wave -position insertpoint  \
sim:/toplevel/Datapat/pre_encoder/din \
sim:/toplevel/Datapat/pre_encoder/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/decoder_block/din \
sim:/toplevel/Datapat/decoder_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/xor_b_mux/sel \
sim:/toplevel/Datapat/xor_b_mux/y
add wave -position insertpoint  \
sim:/toplevel/Datapat/xor_a_mux/sel \
sim:/toplevel/Datapat/xor_a_mux/y
run
run
run
run
run
run -continue
run
run
run
run
restart
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:01
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:11 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 01:33:11 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:11 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 01:33:11 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
vsim work.toplevel
# End time: 03:22:59 on Nov 24,2018, Elapsed time: 0:04:09
# Errors: 0, Warnings: 3
# vsim work.toplevel 
# Start time: 03:22:59 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# WARNING: No extended dataflow license exists
# vsim work.toplevel 
# Start time: 02:21:38 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# vsim work.toplevel 
# Start time: 01:33:56 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# vsim work.toplevel 
# Start time: 01:18:02 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
add wave -position insertpoint  \
sim:/toplevel/FSM_control/ir_data \
sim:/toplevel/FSM_control/next_state \
sim:/toplevel/FSM_control/state
add wave -position insertpoint  \
sim:/toplevel/Datapat/memory_block/memory_block
add wave -position insertpoint  \
sim:/toplevel/Datapat/reg_file_block/registers
add wave -position insertpoint  \
sim:/toplevel/clock \
sim:/toplevel/reset
force -freeze sim:/toplevel/clock 1 0, 0 {50 ps} -r 100
force -freeze sim:/toplevel/reset 1 0
run
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
force -freeze sim:/toplevel/reset 0 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(0) 0110000010000100 0
force -freeze sim:/toplevel/Datapat/reg_file_block/registers(0) 0000000000000100 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(4) 0000000000000001 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(5) 0000000000000111 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(0) 0110000001000001 0
add wave -position insertpoint  \
sim:/toplevel/Datapat/t4_block/din \
sim:/toplevel/Datapat/t4_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/t2_block/din \
sim:/toplevel/Datapat/t2_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/t5_block/din \
sim:/toplevel/Datapat/t5_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/xorblock/dout \
sim:/toplevel/Datapat/xorblock/xor_a \
sim:/toplevel/Datapat/xorblock/xor_b
add wave -position insertpoint  \
sim:/toplevel/Datapat/pre_encoder/din \
sim:/toplevel/Datapat/pre_encoder/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/decoder_block/din \
sim:/toplevel/Datapat/decoder_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/xor_b_mux/sel \
sim:/toplevel/Datapat/xor_b_mux/y
add wave -position insertpoint  \
sim:/toplevel/Datapat/xor_a_mux/sel \
sim:/toplevel/Datapat/xor_a_mux/y
run
run
run
run
run
run -continue
run
run
run
run

# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 02:21:22 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:22 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:01
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 02:21:23 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 02:21:23 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:09 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 01:33:09 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:10 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 01:33:10 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:11 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 01:33:11 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:33:11 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 01:33:11 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
# ERROR: No extended dataflow license exists
# do Datapath_Components_run_msim_rtl_vhdl.do
# if {[file exists rtl_work]} {
# 	vdel -lib rtl_work -all
# }
# vlib rtl_work
# vmap work rtl_work
# Model Technology ModelSim ALTERA vmap 10.4d Lib Mapping Utility 2015.12 Dec 30 2015
# vmap work rtl_work 
# Copying /home/amit/altera_lite/16.0/modelsim_ase/linuxaloem/../modelsim.ini to modelsim.ini
# Modifying modelsim.ini
# 
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TopLevel.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TopLevel
# -- Compiling architecture struct of TopLevel
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/fsm.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package std_logic_arith
# -- Loading package STD_LOGIC_UNSIGNED
# -- Compiling entity fsm
# -- Compiling architecture a1 of fsm
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:56 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg_1b.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg_1b
# -- Compiling architecture struct of reg_1b
# End time: 01:17:56 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/xor.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity xor_block
# -- Compiling architecture Struct of xor_block
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Datapath.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity Datapath
# -- Compiling architecture behave of Datapath
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/alu.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ALU
# -- Compiling architecture ALU_arch of ALU
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1_al.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1_3bit
# -- Compiling architecture Behavioral of mux_4to1_3bit
# -- Compiling entity mux_2to1_3bit
# -- Compiling architecture Behavioral of mux_2to1_3bit
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/TrailZeroes7.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity TrailZeroes7
# -- Compiling architecture Struct of TrailZeroes7
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE9.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE9
# -- Compiling architecture Struct of SE9
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/SE6.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity SE6
# -- Compiling architecture Struct of SE6
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Reg_file.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Reg_file
# -- Compiling architecture behavioral of Reg_file
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Priority_Encoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Priority_Encoder
# -- Compiling architecture priority_enc_arc of Priority_Encoder
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_4to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_4to1
# -- Compiling architecture Behavioral of mux_4to1
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/mux_2to1.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Compiling entity mux_2to1
# -- Compiling architecture Behavioral of mux_2to1
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/memory.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity memory
# -- Compiling architecture struct of memory
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/ir.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity ir
# -- Compiling architecture struct of ir
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/Decoder.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity Decoder
# -- Compiling architecture decoder_arch of Decoder
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# vcom -93 -work work {/home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd}
# Model Technology ModelSim ALTERA vcom 10.4d Compiler 2015.12 Dec 30 2015
# Start time: 01:17:57 on Nov 24,2018
# vcom -reportprogress 300 -93 -work work /home/amit/Desktop/RISC_IITB/Datapath_components/reg.vhd 
# -- Loading package STANDARD
# -- Loading package TEXTIO
# -- Loading package std_logic_1164
# -- Loading package NUMERIC_STD
# -- Compiling entity reg
# -- Compiling architecture struct of reg
# End time: 01:17:57 on Nov 24,2018, Elapsed time: 0:00:00
# Errors: 0, Warnings: 0
# 
# 
# stdin: <EOF>
vsim work.toplevel
# End time: 03:24:08 on Nov 24,2018, Elapsed time: 0:01:09
# Errors: 0, Warnings: 4
# vsim work.toplevel 
# Start time: 03:24:08 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# WARNING: No extended dataflow license exists
# vsim work.toplevel 
# Start time: 02:21:38 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# vsim work.toplevel 
# Start time: 01:33:56 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
# vsim work.toplevel 
# Start time: 01:18:02 on Nov 24,2018
# Loading std.standard
# Loading std.textio(body)
# Loading ieee.std_logic_1164(body)
# Loading work.toplevel(struct)
# Loading work.datapath(behave)
# Loading ieee.numeric_std(body)
# Loading work.decoder(decoder_arch)
# Loading work.priority_encoder(priority_enc_arc)
# Loading work.mux_2to1(behavioral)
# Loading work.memory(struct)
# Loading work.reg(struct)
# Loading work.mux_4to1(behavioral)
# Loading work.reg_1b(struct)
# Loading work.ir(struct)
# Loading work.se6(struct)
# Loading work.se9(struct)
# Loading work.xor_block(struct)
# Loading work.mux_4to1_3bit(behavioral)
# Loading work.reg_file(behavioral)
# Loading work.mux_2to1_3bit(behavioral)
# Loading work.trailzeroes7(struct)
# Loading work.alu(alu_arch)
# Loading ieee.std_logic_arith(body)
# Loading ieee.std_logic_unsigned(body)
# Loading work.fsm(a1)
add wave -position insertpoint  \
sim:/toplevel/FSM_control/ir_data \
sim:/toplevel/FSM_control/next_state \
sim:/toplevel/FSM_control/state
add wave -position insertpoint  \
sim:/toplevel/Datapat/memory_block/memory_block
add wave -position insertpoint  \
sim:/toplevel/Datapat/reg_file_block/registers
add wave -position insertpoint  \
sim:/toplevel/clock \
sim:/toplevel/reset
force -freeze sim:/toplevel/clock 1 0, 0 {50 ps} -r 100
force -freeze sim:/toplevel/reset 1 0
run
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
force -freeze sim:/toplevel/reset 0 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(0) 0110000010000010 0
force -freeze sim:/toplevel/Datapat/reg_file_block/registers(0) 0000000000000100 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(4) 0000000000000001 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(5) 0000000000000111 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(0) 0110000001000001 0
add wave -position insertpoint  \
sim:/toplevel/Datapat/t4_block/din \
sim:/toplevel/Datapat/t4_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/t2_block/din \
sim:/toplevel/Datapat/t2_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/t5_block/din \
sim:/toplevel/Datapat/t5_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/xorblock/dout \
sim:/toplevel/Datapat/xorblock/xor_a \
sim:/toplevel/Datapat/xorblock/xor_b
add wave -position insertpoint  \
sim:/toplevel/Datapat/pre_encoder/din \
sim:/toplevel/Datapat/pre_encoder/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/decoder_block/din \
sim:/toplevel/Datapat/decoder_block/dout
add wave -position insertpoint  \
sim:/toplevel/Datapat/xor_b_mux/sel \
sim:/toplevel/Datapat/xor_b_mux/y
add wave -position insertpoint  \
sim:/toplevel/Datapat/xor_a_mux/sel \
sim:/toplevel/Datapat/xor_a_mux/y
run
run
run
run
run
run -continue
run
run
run
restart
force -freeze sim:/toplevel/clock 1 0, 0 {50 ps} -r 100
force -freeze sim:/toplevel/reset 1 0
run
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/reg_file_block
# ** Warning: NUMERIC_STD.TO_INTEGER: metavalue detected, returning 0
#    Time: 0 ps  Iteration: 0  Instance: /toplevel/Datapat/memory_block
force -freeze sim:/toplevel/reset 0 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(0) 0110000010000010 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(4) 0000000000000011 0
force -freeze sim:/toplevel/Datapat/memory_block/memory_block(5) 0000000000001111 0
force -freeze sim:/toplevel/Datapat/reg_file_block/registers(0) 0000000000000100 0
force -freeze sim:/toplevel/reset 0 0
run
run
run
run
run
run
run
run
run
